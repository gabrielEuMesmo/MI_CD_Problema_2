module N8bits(S,A);

	input [7:0] A;
	output [7:0] S;
	
	not(S[0], A[0]);
	not(S[1], A[1]);
	not(S[2], A[2]);
	not(S[3], A[3]);
	not(S[4], A[4]);
	not(S[5], A[5]);
	not(S[6], A[6]);
	not(S[7], A[7]);
	
endmodule